// list all paths to your design files
`include "../01_RTL/bch.v"
`include "../01_RTL/BMA.v"
`include "../01_RTL/S_calc.v"
