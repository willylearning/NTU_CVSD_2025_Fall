// list all paths to your design files
`include "../01_RTL/IOTDF.v"
`include "../01_RTL/EnDecrypt.v"